`timescale 1ns / 1ps

module mod
#(parameter input_size = 300,
parameter output_size = 256)
    (input clk,
    input reset,
    input [input_size-1:0] x,
    output [output_size-1:0] o);
    
    localparam p44 = 256'd104899928942039473597645237135751317405745389583683433800060134911610808289117;
    localparam p43 = 257'd209799857884078947195290474271502634811490779167366867600120269823221616578234;
    localparam p42 = 258'd419599715768157894390580948543005269622981558334733735200240539646443233156468;
    localparam p41 = 259'd839199431536315788781161897086010539245963116669467470400481079292886466312936;
    localparam p40 = 260'd1678398863072631577562323794172021078491926233338934940800962158585772932625872;
    localparam p39 = 261'd3356797726145263155124647588344042156983852466677869881601924317171545865251744;
    localparam p38 = 262'd6713595452290526310249295176688084313967704933355739763203848634343091730503488;
    localparam p37 = 263'd13427190904581052620498590353376168627935409866711479526407697268686183461006976;
    localparam p36 = 264'd26854381809162105240997180706752337255870819733422959052815394537372366922013952;
    localparam p35 = 265'd53708763618324210481994361413504674511741639466845918105630789074744733844027904;
    localparam p34 = 266'd107417527236648420963988722827009349023483278933691836211261578149489467688055808;
    localparam p33 = 267'd214835054473296841927977445654018698046966557867383672422523156298978935376111616;
    localparam p32 = 268'd429670108946593683855954891308037396093933115734767344845046312597957870752223232;
    localparam p31 = 269'd859340217893187367711909782616074792187866231469534689690092625195915741504446464;
    localparam p30 = 270'd1718680435786374735423819565232149584375732462939069379380185250391831483008892928;
    localparam p29 = 271'd3437360871572749470847639130464299168751464925878138758760370500783662966017785856;
    localparam p28 = 272'd6874721743145498941695278260928598337502929851756277517520741001567325932035571712;
    localparam p27 = 273'd13749443486290997883390556521857196675005859703512555035041482003134651864071143424;
    localparam p26 = 274'd27498886972581995766781113043714393350011719407025110070082964006269303728142286848;
    localparam p25 = 275'd54997773945163991533562226087428786700023438814050220140165928012538607456284573696;
    localparam p24 = 276'd109995547890327983067124452174857573400046877628100440280331856025077214912569147392;
    localparam p23 = 277'd219991095780655966134248904349715146800093755256200880560663712050154429825138294784;
    localparam p22 = 278'd439982191561311932268497808699430293600187510512401761121327424100308859650276589568;
    localparam p21 = 279'd879964383122623864536995617398860587200375021024803522242654848200617719300553179136;
    localparam p20 = 280'd1759928766245247729073991234797721174400750042049607044485309696401235438601106358272;
    localparam p19 = 281'd3519857532490495458147982469595442348801500084099214088970619392802470877202212716544;
    localparam p18 = 282'd7039715064980990916295964939190884697603000168198428177941238785604941754404425433088;
    localparam p17 = 283'd14079430129961981832591929878381769395206000336396856355882477571209883508808850866176;
    localparam p16 = 284'd28158860259923963665183859756763538790412000672793712711764955142419767017617701732352;
    localparam p15 = 285'd56317720519847927330367719513527077580824001345587425423529910284839534035235403464704;
    localparam p14 = 286'd112635441039695854660735439027054155161648002691174850847059820569679068070470806929408;
    localparam p13 = 287'd225270882079391709321470878054108310323296005382349701694119641139358136140941613858816;
    localparam p12 = 288'd450541764158783418642941756108216620646592010764699403388239282278716272281883227717632;
    localparam p11 = 289'd901083528317566837285883512216433241293184021529398806776478564557432544563766455435264;
    localparam p10 = 290'd1802167056635133674571767024432866482586368043058797613552957129114865089127532910870528;
    localparam p9 = 291'd3604334113270267349143534048865732965172736086117595227105914258229730178255065821741056;
    localparam p8 = 292'd7208668226540534698287068097731465930345472172235190454211828516459460356510131643482112;
    localparam p7 = 293'd14417336453081069396574136195462931860690944344470380908423657032918920713020263286964224;
    localparam p6 = 294'd28834672906162138793148272390925863721381888688940761816847314065837841426040526573928448;
    localparam p5 = 295'd57669345812324277586296544781851727442763777377881523633694628131675682852081053147856896;
    localparam p4 = 296'd115338691624648555172593089563703454885527554755763047267389256263351365704162106295713792;
    localparam p3 = 297'd230677383249297110345186179127406909771055109511526094534778512526702731408324212591427584;
    localparam p2 = 298'd461354766498594220690372358254813819542110219023052189069557025053405462816648425182855168;
    localparam p1 = 299'd922709532997188441380744716509627639084220438046104378139114050106810925633296850365710336;
    localparam p0 = 300'd1845419065994376882761489433019255278168440876092208756278228100213621851266593700731420672;
    
    reg [299:0] temp1;
    reg [298:0] temp2;
    reg [297:0] temp3;
    reg [296:0] temp4;
    reg [295:0] temp5;
    reg [294:0] temp6;
    reg [293:0] temp7;
    reg [292:0] temp8;
    reg [291:0] temp9;
    reg [290:0] temp10;
    reg [289:0] temp11;
    reg [288:0] temp12;
    reg [287:0] temp13;
    reg [286:0] temp14;
    reg [285:0] temp15;
    reg [284:0] temp16;
    reg [283:0] temp17;
    reg [282:0] temp18;
    reg [281:0] temp19;
    reg [280:0] temp20;
    reg [279:0] temp21;
    reg [278:0] temp22;
    reg [277:0] temp23;
    reg [276:0] temp24;
    reg [275:0] temp25;
    reg [274:0] temp26;
    reg [273:0] temp27;
    reg [272:0] temp28;
    reg [271:0] temp29;
    reg [270:0] temp30;
    reg [269:0] temp31;
    reg [268:0] temp32;
    reg [267:0] temp33;
    reg [266:0] temp34;
    reg [265:0] temp35;
    reg [264:0] temp36;
    reg [263:0] temp37;
    reg [262:0] temp38;
    reg [261:0] temp39;
    reg [260:0] temp40;
    reg [259:0] temp41;
    reg [258:0] temp42;
    reg [257:0] temp43;
    reg [256:0] temp44;
    reg [255:0] temp_ans;
    
    always@(posedge clk)
        begin
            if(reset == 1)
            begin
                //Flushing the Pipeline
                temp_ans<=0;
                temp1<=0;
                temp2<=0;
                temp3<=0;
                temp4<=0;
                temp5<=0;
                temp6<=0;
                temp7<=0;
                temp8<=0;
                temp9<=0;
                temp10<=0;
                temp11<=0;
                temp12<=0;
                temp13<=0;
                temp14<=0;
                temp15<=0;
                temp16<=0;
                temp17<=0;
                temp18<=0;
                temp19<=0;
                temp20<=0;
                temp21<=0;
                temp22<=0;
                temp23<=0;
                temp24<=0;
                temp25<=0;
                temp26<=0;
                temp27<=0;
                temp28<=0;
                temp29<=0;
                temp30<=0;
                temp31<=0;
                temp32<=0;
                temp33<=0;
                temp34<=0;
                temp35<=0;
                temp36<=0;
                temp37<=0;
                temp38<=0;
                temp39<=0;
                temp40<=0;
                temp41<=0;
                temp42<=0;
                temp43<=0;
                temp44<=0;
            end    
            else
            begin
                temp1<=(x>=p0)?(x-p0):x;
                temp2 <= (temp1>=p1)?(temp1 - p1):temp1;
                temp3 <= (temp2>=p2)?(temp2 - p2):temp2;
                temp4 <= (temp3>=p3)?(temp3 - p3):temp3;
                temp5 <= (temp4>=p4)?(temp4 - p4):temp4;
                temp6 <= (temp5>=p5)?(temp5 - p5):temp5;
                temp7 <= (temp6>=p6)?(temp6 - p6):temp6;
                temp8 <= (temp7>=p7)?(temp7 - p7):temp7;
                temp9 <= (temp8>=p8)?(temp8 - p8):temp8;
                temp10 <= (temp9>=p9)?(temp9 - p9):temp9;
                temp11 <= (temp10>=p10)?(temp10 - p10):temp10;
                temp12 <= (temp11>=p11)?(temp11 - p11):temp11;
                temp13 <= (temp12>=p12)?(temp12 - p12):temp12;
                temp14 <= (temp13>=p13)?(temp13 - p13):temp13;
                temp15 <= (temp14>=p14)?(temp14 - p14):temp14;
                temp16 <= (temp15>=p15)?(temp15 - p15):temp15;
                temp17 <= (temp16>=p16)?(temp16 - p16):temp16;
                temp18 <= (temp17>=p17)?(temp17 - p17):temp17;
                temp19 <= (temp18>=p18)?(temp18 - p18):temp18;
                temp20 <= (temp19>=p19)?(temp19 - p19):temp19;
                temp21 <= (temp20>=p20)?(temp20 - p20):temp20;
                temp22 <= (temp21>=p21)?(temp21 - p21):temp21;
                temp23 <= (temp22>=p22)?(temp22 - p22):temp22;
                temp24 <= (temp23>=p23)?(temp23 - p23):temp23;
                temp25 <= (temp24>=p24)?(temp24 - p24):temp24;
                temp26 <= (temp25>=p25)?(temp25 - p25):temp25;
                temp27 <= (temp26>=p26)?(temp26 - p26):temp26;
                temp28 <= (temp27>=p27)?(temp27 - p27):temp27;
                temp29 <= (temp28>=p28)?(temp28 - p28):temp28;
                temp30 <= (temp29>=p29)?(temp29 - p29):temp29;
                temp31 <= (temp30>=p30)?(temp30 - p30):temp30;
                temp32 <= (temp31>=p31)?(temp31 - p31):temp31;
                temp33 <= (temp32>=p32)?(temp32 - p32):temp32;
                temp34 <= (temp33>=p33)?(temp33 - p33):temp33;
                temp35 <= (temp34>=p34)?(temp34 - p34):temp34;
                temp36 <= (temp35>=p35)?(temp35 - p35):temp35;
                temp37 <= (temp36>=p36)?(temp36 - p36):temp36;
                temp38 <= (temp37>=p37)?(temp37 - p37):temp37;
                temp39 <= (temp38>=p38)?(temp38 - p38):temp38;
                temp40 <= (temp39>=p39)?(temp39 - p39):temp39;
                temp41 <= (temp40>=p40)?(temp40 - p40):temp40;
                temp42 <= (temp41>=p41)?(temp41 - p41):temp41;
                temp43 <= (temp42>=p42)?(temp42 - p42):temp42;
                temp44 <= (temp43>=p43)?(temp43 - p43):temp43;
                temp_ans <= (temp44>=p44)?(temp44 - p44):temp44;
           end     
        end
    assign o = temp_ans;
endmodule

