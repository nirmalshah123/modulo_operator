`timescale 1ns / 1ps

module mod_sims();

    reg clk;
    reg[299:0] inp;
    reg reset = 1'b0;
    wire [255:0] outp;
    
    
    top_level dut(.clk(clk), .reset(reset), .x(inp),.o(outp));
    always #5 clk = ~clk;
    
    initial
        begin
            inp<=0;
            clk = 0;
            #105;
            // Delay of 100 is given, because of GSR(All the FF are at reset for first 100 ns of the start of the device)
            inp<=300'd150524487336639563623712842814162872628549531222968261766193641388199764251004575389192604;
            #10;
            inp<=300'd294959456127685822495157970775287765722667529486654834730625276855868547896099119060820325;
            #10;
            inp<=300'd1202656854464058609431488307863331795492637195567353234051884301400449448732747381894316328;
            #10;
            inp<=300'd1974227788976415422907467170961998261766436360845528330147398301415946167023225814273585185;
            #10;
            inp<=300'd2022472985592125945512641598893286033438697065239165830787352167525645770173646368860661668;
            #10;
            inp<=300'd1023958852955334697519619618737221218739274267451425930995812727592459347644974484832103236;
            #10;
            inp<=300'd1984940186286027590783744038537401932756730753647695780770115433411676647761625635681597594;
            #10;
            inp<=300'd1649871189472749039003995842502815120068594098859429274049633562068646271807712073483709334;
            #10;
            inp<=300'd430489814770949813628430022529264778048747839731404617185964750388739486174008044271307237;
            #10;
            inp<=300'd660615138850469295699441479098126120417373371436076788600343476455587143281957091040534486;
            #10;
            inp<=300'd468882680613132141741494778676518201237710479274385150119175588334468611135133437767129997;
            #10;
            inp<=300'd422612442351370435844979627987617832950830839110997143004225666574390876352949648759508736;
            #10;
            inp<=300'd1189863703862712265048822925171035401497345753236294053482828385621148483886456764009960850;
            #10;
            inp<=300'd991401170101856303843943030205132796264732487024678021386878187077033731984405421162259924;
            #10;
            inp<=300'd1193161160951536389871183986802754472214019327691057865716189468102616654789436589874448705;
            #10;
            inp<=300'd1580228807310313234863430114426460376313011936423405452812905023475779144570326695994909710;
            #10;
            inp<=300'd1228810452864306047510288545604077269082868803300272191858981428676649298973334928189395747;
            #10;
            inp<=300'd446418310676693138243630173800033054437830559031403991152639861006386416091703402950158073;
            #10;
            inp<=300'd2022878969739416693936904418302648811821431057329484800244786472173690680244182877283461312;
            #10;
            inp<=300'd1916085352928700927882483843489998815220091427491777183225691145293478331240686981477707149;
            #10;
            inp<=300'd1610755061310521337308566166725900057304787515566021868235378878999821126599418101176254234;
            #10;
            inp<=300'd1336379611678207369486583950548099693629148595966744723016742452348707848714414350190086289;
            #10;
            inp<=300'd1507123749315590798000268541694215572584570265631236368511750394964111993762630945066422477;
            #10;
            inp<=300'd206954447307206413370152646333148319446437416468990496630445900066391040141111002655710855;
            #10;
            inp<=300'd236266677382387956749660761470674459152862745698863372073314140313501109847676698194129595;
            #10;
            inp<=300'd1276200268074128046154313081829850013593125970511160765957460806455894275504275504148581388;
            #10;
            inp<=300'd1279595098809861645268276665467561517377484732584479603520310638150355730912251819976717319;
            #10;
            inp<=300'd416536838574030759825757340526186725887375246092638814792655306682035377770952730181264637;
            #10;
            inp<=300'd2021679642816327682571435047790229735552101977319087831472411933541610950718649498930905053;
            #10;
            inp<=300'd885980994237117076908327713215529478739446202197784648456231279145190506761054294943792769;
            #10;
            inp<=300'd740612501472875269447729741320127863544213181809872739021537004510497588853111872585447210;
            #10;
            inp<=300'd113309578167685667991561476704339694238816997238889357596725876542163739955021957268293743;
            #10;
            inp<=300'd667970426667450325978309081261230951982458738169454009042067661551363104993042199433345027;
            #10;
            inp<=300'd633675655809992050254798722050815608305170676100678295742096533026983846108988884224430677;
            #10;
            inp<=300'd892468545387626262968691877775941926452467634001594648906758492620732180283989195767456032;
            #10;
            inp<=300'd858693702366366517340345752701860622914237011630118417149404381625403441290378876439961400;
            #10;
            inp<=300'd915585280745245623231501888061240230077914864677901661196143916074112433211000025810267743;
            #10;
            inp<=300'd1926646893752414275441407664434711233710683383684690336585035824889588598243013353138717624;
            #10;
            inp<=300'd665967352423373847357036400525633876105906116114946906936860344013829639622331140033805907;
            #10;
            inp<=300'd1846839987257100878514842443983592805839232265680020647729645918379729209321610001823119550;
            #10;
            
        # 100000;
            $finish;
        end
endmodule
//Input in hex is
//0x12eab58c2946605e6db09a51f84c0e5b11b6c52fcebb8bdfab7afc8f50cb1ab61cba1e2119c
//0x25118142585ae00d9f035e36baa3bdff1f5951f343a0c1aa08644a3c879c413f20543552165
//0x972428ab8234c7f3d97c64f8f7b4c4289306cae4875184536df7754e59479e6f2384d888128
//0xf81b51fb487bfed6162f447522575732c5a5d1b8b36bc5dc8638f07a2633bec04866de17021
//0xfe2b79ddca2b2a64763f11bc62802caa7203834327fbfe9dfa4ba7bfb40c99f259fbd61e7a4
//0x80af0b76b73701005fdf8b7cefb1a0fe852e387ed7424adb8b12288b6766d9b2c26a707ab44
//0xf973f645dc2b35da5c0f71bc3ff7c245d404aae75c57f46cd35dfa610b5155d681b89ddf89a
//0xcf580b240d0d2e10c9858f1e20ca9a4fe465d22a130a442dbd18600d07f3363a4ee43666b96
//0x3619d1c7f8d4f0ab6bbb54637226d6f2d837a353486b6d2b3cfa47cec2f9e08f521169209e5
//0x530577279c7c5f8cff8e452819d227cd5d2826e2f363bcb7f62dd05b16635b484af3e1b9fd6
//0x3aed00f63c385fbafdd240ba3323d2e3a372f00aff8ee277abafc1c75941d6f643d798f1b8d
//0x351c63041ba91b0143a4f701daa7d7a18c83ed3b5c6acc9bba30fa4943aadad8cc4a5d8cf00
//0x9588931a5135d2aa91f3f75088bb0168b33b654712719b155f0f829e6d4c45676e7eaba5592
//0x7c97976345d7d7542b10a2c4d3ba2c5977a02494097cc3da33feac6ba520365dac6e58465d4
//0x95f2a943629a3de1e6fd857b1ba36adad2204e648fb658fadce9a656568f53466fa30a18941
//0xc6977e1073bb9b4113aebfa53656b4fe2738998bf705a45aceb91afde7d270ac73d24d2e40e
//0x9a6d941dc2e15886229c4d012461fcc01b3c81a7d771249f10a44246cab24293324543d9323
//0x381a465753c709acbcea8d027956c547c3e2ad06615c1dc00355df78b0ba3d29e8bd349e6f9
//0xfe388996d6965a49774e236ff73ddc964021885eef19b7b2cec533672ab6e349b313696a8c0
//0xf0ccbf8556fe358cd05710fa87a394389570205bad4fd52d1799058f95e8c5495c55b162d8d
//0xca6d971ae11260c1c046dad06f79ff8821e51f753f41a498f488a57230ecaa58c9921e4bf1a
//0xa7f2519eb8ca8bd11104f9e3718aff4982915a256fd35fc3ac029392a933b2052f748a58891
//0xbd678a120bb5906b9615b2018604fbb3974f947a196003c86d1ec68716ec3d63b4275ab90cd
//0x1a022fe5bfb72395488c6c3771924be7993f1d5a81177fb9d315c9ee8eaa66c112f23315e87
//0x1db13a201226c361d6e18c11ccc1a77e300c5fb1ae5914978f430158de6ec4ae7f76df0b2bb
//0xa06237003f8e2a2db01e918a867a00a36bf8aba0d76930855192c17d5d91d75361b0fe10c0c
//0xa0cf6f23c4ab2296b88385597e9cf694358ccee34fe50130886c065d37ee5dcc3117c727407
//0x3458ebc89437ec25dad7be658fe8a815572a1de44610d28f6e1de168fd45d9c6d11513664fd
//0xfe11f3d2794f0033b648ae290296d6bb17df74dcf9f6c1eab10594d89b62fc9f0309121ffdd
//0x6f57fd1b099e7219b5884634f3c10e66ec0fc0a9739fd61a31db8ed98ecb7ead0763850fe81
//0x5d1328cdf39e22a48a791eba18384a16814dc824a0ad327476d5a3e04808a431c40b36fb72a
//0xe3d6c2061ac8704f0aab19473e1fa021d6a1c23551c6a08d5d0025b1ff3b1db005f738c86f
//0x53f219fba16744416c20f4407cf36989887a61be15feae1610d83bee96f3fd7c66874b27803
//0x4fa2c3171231a8967c7cb1ca94aa4006d235203a953c79a958c4c981896379115827781d255
//0x7028b52cb777f405bbd5f717b9e5b8c8ee4b09d600234fcd64c9907d6c6b98c29d2cd94a120
//0x6bea18749720ae899b6f0b0196be9b464d5de856b040272d48791d113ce0f76795fde9f1f38
//0x73106cbcb4768c995eb7680cee30ef9178e0a092402dc5ca6de2e829073cbc474c7c228ee5f
//0xf2208958212fcd10fdce97fc85fa8ac685d870c14777f0c6b248d22defb3116b99f619a83b8
//0x53b1a87a9863dc624a0831b905d085d92c8aade74fff65df0cbb2f3187ade182c18921cfe53
//0xe818f84f070cca6ac732160541671f4ae14850aada15283dd4395d40929536f880ce42538be




//Answers are
//0xd9c30588b3715290d80fbe34b447b83ca4be1dbf1d976b59f0d7bfb70a246c60
//0x144425fe7b7bebbcfa54c3ea5dd3c2c9f3df066f0caf1fe253ed1dbbd617d038
//0x8227c5b47211d03dc6c41bb2cd2e65e001f2981d24322c7f508624eb2568562e
//0xf92c95cd512629f1fcfe5768aab9c48ed7da6a7ebee9f5a5104e5e35b49853e
//0x2ac3a83514c8f1a2e08f95ebcc9968d3977e3a442869dde781a660b1a6d04d90
//0xb782df2b07d44e83f73f104655fc860944ced6ec045ca2cba2e319c6f358954c
//0x71ff55c6226f7ea52ca716baa48251acec7176433dc3e8ce646877070ee5239d
//0x16425df805bc6b3cb4bff525268870139e9b308b2dfec543104380fd0d8e7d16
//0x144a010089bf688596d9373115b3afa0c4802c44da7804f04d3130f93122b87e
//0x742fb03f59b8cb2df21bfbc6a190b09fda12156997a99abe1aef94de383184b4
//0xb36512b5f7ba8ce1645578e40614a54c17f62db26aad63e9478dd4dbe7a63eed
//0x73d3ee122e342a8e498433047aa257948e3c94ef421a37749f7cf3502d463e34
//0x837e18739ae0c267306484135592df0759ac9d73fa03da777a44051a4bcadc4
//0xe11d8fee13e15e366aa39c8be6adaaa9416012ad6e3dcad4b33f1d418fe649bc
//0xbb912b4ce07587bdd189590a982a8e84d9c45ed276642be6ac0bc7b4183cc65c
//0x28c658c7c46b95d63ecce81b37dad7f402484e1c926f3f48ee0e046456fae969
//0xbfdcf12cc1ff7892a470d5d7f7cdcdc2f0346d36511f5a501a15282f2c3d646e
//0xa613d52dd827a93e03cc6022069f85d38f606d54962826cb0f04c2f9a6784d85
//0x85c74264652bcc25db84c89caa91c8d6ffbd75e8fc1471eda4e082323ce9f554
//0x2307b7339e34ff8d2b6427770dbdb0b8c0a7c5bd2c73c7db22fc23f2d843961d
//0xcea10ce08cb4b6d605c3831d6240c3b50b5ef40ca4ced7fcf65cc3d31865d0d7
//0xab218d7872b6b264bc756bc89d271142aba8a578eefb6faf8cc4bccea95c4e3b
//0xb93afa7e12b4a7b415a2058ce34fe7a9bebf7d80fa3f598ffebe51d3a2e9322c
//0xbe51c475e6a9a5d3c0a19cf435e86bfd4305b5e4ad527a6b7f90aab77df3f609
//0x96d210b8940d5444443c029d41ba782023cf74218dc66d0e8798127c76c4a7b5
//0xba5e0cf4d45738f49f38a47ebf12958155a413d83b94b84618000b84498db837
//0xba052bb28cc95afa428507e406a5526f67d69dd3df57436e89d55ec338c01496
//0x4fcaace4fd0452838ecba2fe9f6d8164f1452d9bd3128131ed360bda7a80783e
//0xc2e18e40a05a7de244d870c1dfcf60277ae45beed985762ddb0067c444975571
//0x75153455bc1f68af57b899e3517d496125058f47cc23c10d452d39a1ce495fc
//0x8f03dcae06974c71b18ac997f1c6f880d09e05a0047fa9bd2ae9aabd3be9244e
//0x8a897bdd5e45e3efd5dde146f97710f598b1dc24b8177e0399d9f8c98f2908bb
//0xb3c3a3e6a5dfdb83fbfef473d926ef1fd94cfefeeb4da718a550f2c7b4d49b18
//0x876c33685429414bd3db218d1e851926f07c1af26f5b3698b3d767fbbd8a783b
//0x41582055634dcef7e4345cbb95140378d82a64b89ac1c60d68e5ad95c3cfae78
//0xda87aa51a5aeeccf4fce4d062cea8602a95112b3bd0182eea5b092a6567e8d40
//0x933901539fbea6671c5a9458b4febac26c86d1919c92a794a9072c0d95ea7c34
//0x16e6d7ec158ddc9379876fc2f8db17912536b2ec0f8c42704f4ef2baa06dbab2
//0x9f7993c4832d4922d2b55fcbf0b21daef27a8a31d9ae01e895e61960e49fe7df
//0xd8e7c19cbf16c0605bb1793b97f624d005e03ab648511313469677173b719d24


