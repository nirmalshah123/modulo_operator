`timescale 1ns / 1ps

module mac(
    input clk,
    input[299:0] x,
    output[260:0] o,
    input reset
    );
    localparam x0 = 1'd1;
    localparam x1 = 2'd2;
    localparam x2 = 3'd4;
    localparam x3 = 4'd8;
    localparam x4 = 5'd16;
    localparam x5 = 6'd32;
    localparam x6 = 7'd64;
    localparam x7 = 8'd128;
    localparam x8 = 9'd256;
    localparam x9 = 10'd512;
    localparam x10 = 11'd1024;
    localparam x11 = 12'd2048;
    localparam x12 = 13'd4096;
    localparam x13 = 14'd8192;
    localparam x14 = 15'd16384;
    localparam x15 = 16'd32768;
    localparam x16 = 17'd65536;
    localparam x17 = 18'd131072;
    localparam x18 = 19'd262144;
    localparam x19 = 20'd524288;
    localparam x20 = 21'd1048576;
    localparam x21 = 22'd2097152;
    localparam x22 = 23'd4194304;
    localparam x23 = 24'd8388608;
    localparam x24 = 25'd16777216;
    localparam x25 = 26'd33554432;
    localparam x26 = 27'd67108864;
    localparam x27 = 28'd134217728;
    localparam x28 = 29'd268435456;
    localparam x29 = 30'd536870912;
    localparam x30 = 31'd1073741824;
    localparam x31 = 32'd2147483648;
    localparam x32 = 33'd4294967296;
    localparam x33 = 34'd8589934592;
    localparam x34 = 35'd17179869184;
    localparam x35 = 36'd34359738368;
    localparam x36 = 37'd68719476736;
    localparam x37 = 38'd137438953472;
    localparam x38 = 39'd274877906944;
    localparam x39 = 40'd549755813888;
    localparam x40 = 41'd1099511627776;
    localparam x41 = 42'd2199023255552;
    localparam x42 = 43'd4398046511104;
    localparam x43 = 44'd8796093022208;
    localparam x44 = 45'd17592186044416;
    localparam x45 = 46'd35184372088832;
    localparam x46 = 47'd70368744177664;
    localparam x47 = 48'd140737488355328;
    localparam x48 = 49'd281474976710656;
    localparam x49 = 50'd562949953421312;
    localparam x50 = 51'd1125899906842624;
    localparam x51 = 52'd2251799813685248;
    localparam x52 = 53'd4503599627370496;
    localparam x53 = 54'd9007199254740992;
    localparam x54 = 55'd18014398509481984;
    localparam x55 = 56'd36028797018963968;
    localparam x56 = 57'd72057594037927936;
    localparam x57 = 58'd144115188075855872;
    localparam x58 = 59'd288230376151711744;
    localparam x59 = 60'd576460752303423488;
    localparam x60 = 61'd1152921504606846976;
    localparam x61 = 62'd2305843009213693952;
    localparam x62 = 63'd4611686018427387904;
    localparam x63 = 64'd9223372036854775808;
    localparam x64 = 65'd18446744073709551616;
    localparam x65 = 66'd36893488147419103232;
    localparam x66 = 67'd73786976294838206464;
    localparam x67 = 68'd147573952589676412928;
    localparam x68 = 69'd295147905179352825856;
    localparam x69 = 70'd590295810358705651712;
    localparam x70 = 71'd1180591620717411303424;
    localparam x71 = 72'd2361183241434822606848;
    localparam x72 = 73'd4722366482869645213696;
    localparam x73 = 74'd9444732965739290427392;
    localparam x74 = 75'd18889465931478580854784;
    localparam x75 = 76'd37778931862957161709568;
    localparam x76 = 77'd75557863725914323419136;
    localparam x77 = 78'd151115727451828646838272;
    localparam x78 = 79'd302231454903657293676544;
    localparam x79 = 80'd604462909807314587353088;
    localparam x80 = 81'd1208925819614629174706176;
    localparam x81 = 82'd2417851639229258349412352;
    localparam x82 = 83'd4835703278458516698824704;
    localparam x83 = 84'd9671406556917033397649408;
    localparam x84 = 85'd19342813113834066795298816;
    localparam x85 = 86'd38685626227668133590597632;
    localparam x86 = 87'd77371252455336267181195264;
    localparam x87 = 88'd154742504910672534362390528;
    localparam x88 = 89'd309485009821345068724781056;
    localparam x89 = 90'd618970019642690137449562112;
    localparam x90 = 91'd1237940039285380274899124224;
    localparam x91 = 92'd2475880078570760549798248448;
    localparam x92 = 93'd4951760157141521099596496896;
    localparam x93 = 94'd9903520314283042199192993792;
    localparam x94 = 95'd19807040628566084398385987584;
    localparam x95 = 96'd39614081257132168796771975168;
    localparam x96 = 97'd79228162514264337593543950336;
    localparam x97 = 98'd158456325028528675187087900672;
    localparam x98 = 99'd316912650057057350374175801344;
    localparam x99 = 100'd633825300114114700748351602688;
    localparam x100 = 101'd1267650600228229401496703205376;
    localparam x101 = 102'd2535301200456458802993406410752;
    localparam x102 = 103'd5070602400912917605986812821504;
    localparam x103 = 104'd10141204801825835211973625643008;
    localparam x104 = 105'd20282409603651670423947251286016;
    localparam x105 = 106'd40564819207303340847894502572032;
    localparam x106 = 107'd81129638414606681695789005144064;
    localparam x107 = 108'd162259276829213363391578010288128;
    localparam x108 = 109'd324518553658426726783156020576256;
    localparam x109 = 110'd649037107316853453566312041152512;
    localparam x110 = 111'd1298074214633706907132624082305024;
    localparam x111 = 112'd2596148429267413814265248164610048;
    localparam x112 = 113'd5192296858534827628530496329220096;
    localparam x113 = 114'd10384593717069655257060992658440192;
    localparam x114 = 115'd20769187434139310514121985316880384;
    localparam x115 = 116'd41538374868278621028243970633760768;
    localparam x116 = 117'd83076749736557242056487941267521536;
    localparam x117 = 118'd166153499473114484112975882535043072;
    localparam x118 = 119'd332306998946228968225951765070086144;
    localparam x119 = 120'd664613997892457936451903530140172288;
    localparam x120 = 121'd1329227995784915872903807060280344576;
    localparam x121 = 122'd2658455991569831745807614120560689152;
    localparam x122 = 123'd5316911983139663491615228241121378304;
    localparam x123 = 124'd10633823966279326983230456482242756608;
    localparam x124 = 125'd21267647932558653966460912964485513216;
    localparam x125 = 126'd42535295865117307932921825928971026432;
    localparam x126 = 127'd85070591730234615865843651857942052864;
    localparam x127 = 128'd170141183460469231731687303715884105728;
    localparam x128 = 129'd340282366920938463463374607431768211456;
    localparam x129 = 130'd680564733841876926926749214863536422912;
    localparam x130 = 131'd1361129467683753853853498429727072845824;
    localparam x131 = 132'd2722258935367507707706996859454145691648;
    localparam x132 = 133'd5444517870735015415413993718908291383296;
    localparam x133 = 134'd10889035741470030830827987437816582766592;
    localparam x134 = 135'd21778071482940061661655974875633165533184;
    localparam x135 = 136'd43556142965880123323311949751266331066368;
    localparam x136 = 137'd87112285931760246646623899502532662132736;
    localparam x137 = 138'd174224571863520493293247799005065324265472;
    localparam x138 = 139'd348449143727040986586495598010130648530944;
    localparam x139 = 140'd696898287454081973172991196020261297061888;
    localparam x140 = 141'd1393796574908163946345982392040522594123776;
    localparam x141 = 142'd2787593149816327892691964784081045188247552;
    localparam x142 = 143'd5575186299632655785383929568162090376495104;
    localparam x143 = 144'd11150372599265311570767859136324180752990208;
    localparam x144 = 145'd22300745198530623141535718272648361505980416;
    localparam x145 = 146'd44601490397061246283071436545296723011960832;
    localparam x146 = 147'd89202980794122492566142873090593446023921664;
    localparam x147 = 148'd178405961588244985132285746181186892047843328;
    localparam x148 = 149'd356811923176489970264571492362373784095686656;
    localparam x149 = 150'd713623846352979940529142984724747568191373312;
    localparam x150 = 151'd1427247692705959881058285969449495136382746624;
    localparam x151 = 152'd2854495385411919762116571938898990272765493248;
    localparam x152 = 153'd5708990770823839524233143877797980545530986496;
    localparam x153 = 154'd11417981541647679048466287755595961091061972992;
    localparam x154 = 155'd22835963083295358096932575511191922182123945984;
    localparam x155 = 156'd45671926166590716193865151022383844364247891968;
    localparam x156 = 157'd91343852333181432387730302044767688728495783936;
    localparam x157 = 158'd182687704666362864775460604089535377456991567872;
    localparam x158 = 159'd365375409332725729550921208179070754913983135744;
    localparam x159 = 160'd730750818665451459101842416358141509827966271488;
    localparam x160 = 161'd1461501637330902918203684832716283019655932542976;
    localparam x161 = 162'd2923003274661805836407369665432566039311865085952;
    localparam x162 = 163'd5846006549323611672814739330865132078623730171904;
    localparam x163 = 164'd11692013098647223345629478661730264157247460343808;
    localparam x164 = 165'd23384026197294446691258957323460528314494920687616;
    localparam x165 = 166'd46768052394588893382517914646921056628989841375232;
    localparam x166 = 167'd93536104789177786765035829293842113257979682750464;
    localparam x167 = 168'd187072209578355573530071658587684226515959365500928;
    localparam x168 = 169'd374144419156711147060143317175368453031918731001856;
    localparam x169 = 170'd748288838313422294120286634350736906063837462003712;
    localparam x170 = 171'd1496577676626844588240573268701473812127674924007424;
    localparam x171 = 172'd2993155353253689176481146537402947624255349848014848;
    localparam x172 = 173'd5986310706507378352962293074805895248510699696029696;
    localparam x173 = 174'd11972621413014756705924586149611790497021399392059392;
    localparam x174 = 175'd23945242826029513411849172299223580994042798784118784;
    localparam x175 = 176'd47890485652059026823698344598447161988085597568237568;
    localparam x176 = 177'd95780971304118053647396689196894323976171195136475136;
    localparam x177 = 178'd191561942608236107294793378393788647952342390272950272;
    localparam x178 = 179'd383123885216472214589586756787577295904684780545900544;
    localparam x179 = 180'd766247770432944429179173513575154591809369561091801088;
    localparam x180 = 181'd1532495540865888858358347027150309183618739122183602176;
    localparam x181 = 182'd3064991081731777716716694054300618367237478244367204352;
    localparam x182 = 183'd6129982163463555433433388108601236734474956488734408704;
    localparam x183 = 184'd12259964326927110866866776217202473468949912977468817408;
    localparam x184 = 185'd24519928653854221733733552434404946937899825954937634816;
    localparam x185 = 186'd49039857307708443467467104868809893875799651909875269632;
    localparam x186 = 187'd98079714615416886934934209737619787751599303819750539264;
    localparam x187 = 188'd196159429230833773869868419475239575503198607639501078528;
    localparam x188 = 189'd392318858461667547739736838950479151006397215279002157056;
    localparam x189 = 190'd784637716923335095479473677900958302012794430558004314112;
    localparam x190 = 191'd1569275433846670190958947355801916604025588861116008628224;
    localparam x191 = 192'd3138550867693340381917894711603833208051177722232017256448;
    localparam x192 = 193'd6277101735386680763835789423207666416102355444464034512896;
    localparam x193 = 194'd12554203470773361527671578846415332832204710888928069025792;
    localparam x194 = 195'd25108406941546723055343157692830665664409421777856138051584;
    localparam x195 = 196'd50216813883093446110686315385661331328818843555712276103168;
    localparam x196 = 197'd100433627766186892221372630771322662657637687111424552206336;
    localparam x197 = 198'd200867255532373784442745261542645325315275374222849104412672;
    localparam x198 = 199'd401734511064747568885490523085290650630550748445698208825344;
    localparam x199 = 200'd803469022129495137770981046170581301261101496891396417650688;
    localparam x200 = 201'd1606938044258990275541962092341162602522202993782792835301376;
    localparam x201 = 202'd3213876088517980551083924184682325205044405987565585670602752;
    localparam x202 = 203'd6427752177035961102167848369364650410088811975131171341205504;
    localparam x203 = 204'd12855504354071922204335696738729300820177623950262342682411008;
    localparam x204 = 205'd25711008708143844408671393477458601640355247900524685364822016;
    localparam x205 = 206'd51422017416287688817342786954917203280710495801049370729644032;
    localparam x206 = 207'd102844034832575377634685573909834406561420991602098741459288064;
    localparam x207 = 208'd205688069665150755269371147819668813122841983204197482918576128;
    localparam x208 = 209'd411376139330301510538742295639337626245683966408394965837152256;
    localparam x209 = 210'd822752278660603021077484591278675252491367932816789931674304512;
    localparam x210 = 211'd1645504557321206042154969182557350504982735865633579863348609024;
    localparam x211 = 212'd3291009114642412084309938365114701009965471731267159726697218048;
    localparam x212 = 213'd6582018229284824168619876730229402019930943462534319453394436096;
    localparam x213 = 214'd13164036458569648337239753460458804039861886925068638906788872192;
    localparam x214 = 215'd26328072917139296674479506920917608079723773850137277813577744384;
    localparam x215 = 216'd52656145834278593348959013841835216159447547700274555627155488768;
    localparam x216 = 217'd105312291668557186697918027683670432318895095400549111254310977536;
    localparam x217 = 218'd210624583337114373395836055367340864637790190801098222508621955072;
    localparam x218 = 219'd421249166674228746791672110734681729275580381602196445017243910144;
    localparam x219 = 220'd842498333348457493583344221469363458551160763204392890034487820288;
    localparam x220 = 221'd1684996666696914987166688442938726917102321526408785780068975640576;
    localparam x221 = 222'd3369993333393829974333376885877453834204643052817571560137951281152;
    localparam x222 = 223'd6739986666787659948666753771754907668409286105635143120275902562304;
    localparam x223 = 224'd13479973333575319897333507543509815336818572211270286240551805124608;
    localparam x224 = 225'd26959946667150639794667015087019630673637144422540572481103610249216;
    localparam x225 = 226'd53919893334301279589334030174039261347274288845081144962207220498432;
    localparam x226 = 227'd107839786668602559178668060348078522694548577690162289924414440996864;
    localparam x227 = 228'd215679573337205118357336120696157045389097155380324579848828881993728;
    localparam x228 = 229'd431359146674410236714672241392314090778194310760649159697657763987456;
    localparam x229 = 230'd862718293348820473429344482784628181556388621521298319395315527974912;
    localparam x230 = 231'd1725436586697640946858688965569256363112777243042596638790631055949824;
    localparam x231 = 232'd3450873173395281893717377931138512726225554486085193277581262111899648;
    localparam x232 = 233'd6901746346790563787434755862277025452451108972170386555162524223799296;
    localparam x233 = 234'd13803492693581127574869511724554050904902217944340773110325048447598592;
    localparam x234 = 235'd27606985387162255149739023449108101809804435888681546220650096895197184;
    localparam x235 = 236'd55213970774324510299478046898216203619608871777363092441300193790394368;
    localparam x236 = 237'd110427941548649020598956093796432407239217743554726184882600387580788736;
    localparam x237 = 238'd220855883097298041197912187592864814478435487109452369765200775161577472;
    localparam x238 = 239'd441711766194596082395824375185729628956870974218904739530401550323154944;
    localparam x239 = 240'd883423532389192164791648750371459257913741948437809479060803100646309888;
    localparam x240 = 241'd1766847064778384329583297500742918515827483896875618958121606201292619776;
    localparam x241 = 242'd3533694129556768659166595001485837031654967793751237916243212402585239552;
    localparam x242 = 243'd7067388259113537318333190002971674063309935587502475832486424805170479104;
    localparam x243 = 244'd14134776518227074636666380005943348126619871175004951664972849610340958208;
    localparam x244 = 245'd28269553036454149273332760011886696253239742350009903329945699220681916416;
    localparam x245 = 246'd56539106072908298546665520023773392506479484700019806659891398441363832832;
    localparam x246 = 247'd113078212145816597093331040047546785012958969400039613319782796882727665664;
    localparam x247 = 248'd226156424291633194186662080095093570025917938800079226639565593765455331328;
    localparam x248 = 249'd452312848583266388373324160190187140051835877600158453279131187530910662656;
    localparam x249 = 250'd904625697166532776746648320380374280103671755200316906558262375061821325312;
    localparam x250 = 251'd1809251394333065553493296640760748560207343510400633813116524750123642650624;
    localparam x251 = 252'd3618502788666131106986593281521497120414687020801267626233049500247285301248;
    localparam x252 = 253'd7237005577332262213973186563042994240829374041602535252466099000494570602496;
    localparam x253 = 254'd14474011154664524427946373126085988481658748083205070504932198000989141204992;
    localparam x254 = 255'd28948022309329048855892746252171976963317496166410141009864396001978282409984;
    localparam x255 = 256'd57896044618658097711785492504343953926634992332820282019728792003956564819968;
    localparam x256 = 253'd10892160295276721825925747872936590447524595081957130239397449096302321350819;
    localparam x257 = 254'd21784320590553443651851495745873180895049190163914260478794898192604642701638;
    localparam x258 = 255'd43568641181106887303702991491746361790098380327828520957589796385209285403276;
    localparam x259 = 256'd87137282362213774607405982983492723580196760655657041915179592770418570806552;
    localparam x260 = 256'd69374635782388075617166728831234129754648131727630650030299050629226333323987;
    localparam x261 = 255'd33849342622736677636688220526716942103550873871577866260537966346841858358857;
    localparam x262 = 256'd67698685245473355273376441053433884207101747743155732521075932693683716717714;
    localparam x263 = 255'd30497441548907236949107644971116451008458105902628031242091730475756625146311;
    localparam x264 = 256'd60994883097814473898215289942232902016916211805256062484183460951513250292622;
    localparam x265 = 254'd17089837253589474198785342748714486628087034026828691168306786991415692296127;
    localparam x266 = 255'd34179674507178948397570685497428973256174068053657382336613573982831384592254;
    localparam x267 = 256'd68359349014357896795141370994857946512348136107314764673227147965662769184508;
    localparam x268 = 255'd31818769086676319992637504853964575618950882630946095546394161019714730079899;
    localparam x269 = 256'd63637538173352639985275009707929151237901765261892191092788322039429460159798;
    localparam x270 = 254'd22375147404665806372904782280106985070058140940100948385516509167248112030479;
    localparam x271 = 255'd44750294809331612745809564560213970140116281880201896771033018334496224060958;
    localparam x272 = 256'd89500589618663225491619129120427940280232563760403793542066036668992448121916;
    localparam x273 = 256'd74101250295286977385593021105104563154719737937124153284071938426374087954715;
    localparam x274 = 255'd43302571648534481173540805074457808903694086290564872768083741941137367620313;
    localparam x275 = 256'd86605143297068962347081610148915617807388172581129745536167483882274735240626;
    localparam x276 = 256'd68310357652098451096517983162079918209030955578576057272274832852938662192135;
    localparam x277 = 255'd31720786362157428595390729188408519012316521573468680744489530794266516095153;
    localparam x278 = 256'd63441572724314857190781458376817038024633043146937361488979061588533032190306;
    localparam x279 = 254'd21983216506590240783917679617882758643520696710191289177897988265455256091495;
    localparam x280 = 255'd43966433013180481567835359235765517287041393420382578355795976530910512182990;
    localparam x281 = 256'd87932866026360963135670718471531034574082786840765156711591953061821024365980;
    localparam x282 = 256'd70965803110682452673696199807310751742420184097846879623123771212031240442843;
    localparam x283 = 255'd37031677279325431749747162478870186079094978612010325446187407512451672596569;
    localparam x284 = 256'd74063354558650863499494324957740372158189957224020650892374815024903345193138;
    localparam x285 = 255'd43226780175262253401343412779729426910634524864357867984689495138195882097159;
    localparam x286 = 256'd86453560350524506802686825559458853821269049728715735969378990276391764194318;
    localparam x287 = 256'd68007191759009540007728413983166390236792709873748038138697845641172720099519;
    localparam x288 = 255'd31114454575979606417811590830581463067840030163812642477335556370734631909921;
    localparam x289 = 256'd62228909151959212835623181661162926135680060327625284954671112741469263819842;
    localparam x290 = 254'd19557889361878952073601126186574534865614731071567136109282090571327719350567;
    localparam x291 = 255'd39115778723757904147202252373149069731229462143134272218564181142655438701134;
    localparam x292 = 256'd78231557447515808294404504746298139462458924286268544437128362285310877402268;
    localparam x293 = 255'd51563185952992142991163772356844961519172458988853655074196589659010946515419;
    localparam x294 = 256'd103126371905984285982327544713689923038344917977707310148393179318021893030838;
    localparam x295 = 256'd101352814869929098367009852291628528670944446371731186496726223724432977772559;
    localparam x296 = 256'd97805700797818723136374467447505739936143503159778939193392312537255147256001;
    localparam x297 = 256'd90711472653597972675103697759260162466541616735874444586724490162899486222885;
    localparam x298 = 256'd76523016365156471752562158382769007527337843888065455373388845414188164156653;
    localparam x299 = 255'd48146103788273469907479079629786697648930298192447476946717555916765520024189;

    
    reg [260:0] temp0 = 0;
    reg [260:0] temp1 = 0;
    reg [260:0] temp2 = 0;
    reg [260:0] temp3 = 0;
    reg [260:0] temp4 = 0;
    reg [260:0] temp5 = 0;
    reg [260:0] temp6 = 0;
    reg [260:0] temp7 = 0;
    reg [260:0] temp8 = 0;
    reg [260:0] temp9 = 0;
    reg [260:0] temp10 = 0;
    reg [260:0] temp11 = 0;
    reg [260:0] temp12 = 0;
    reg [260:0] temp13 = 0;
    reg [260:0] temp14 = 0;
    reg [260:0] temp15 = 0;
    reg [260:0] temp16 = 0;
    reg [260:0] temp17 = 0;
    reg [260:0] temp18 = 0;
    reg [260:0] temp19 = 0;
    reg [260:0] temp20 = 0;
    reg [260:0] temp21 = 0;
    reg [260:0] temp22 = 0;
    reg [260:0] temp23 = 0;
    reg [260:0] temp24 = 0;
    reg [260:0] temp25 = 0;
    reg [260:0] temp26 = 0;
    reg [260:0] temp27 = 0;
    reg [260:0] temp28 = 0;
    reg [260:0] temp29 = 0;
    reg [260:0] temp30 = 0;
    reg [260:0] temp31 = 0;
    reg [260:0] temp32 = 0;
    reg [260:0] temp33 = 0;
    reg [260:0] temp34 = 0;
    reg [260:0] temp35 = 0;
    reg [260:0] temp36 = 0;
    reg [260:0] temp37 = 0;
    reg [260:0] temp38 = 0;
    reg [260:0] temp39 = 0;
    reg [260:0] temp40 = 0;
    reg [260:0] temp41 = 0;
    reg [260:0] temp42 = 0;
    reg [260:0] temp43 = 0;
    reg [260:0] temp44 = 0;
    reg [260:0] temp45 = 0;
    reg [260:0] temp46 = 0;
    reg [260:0] temp47 = 0;
    reg [260:0] temp48 = 0;
    reg [260:0] temp49 = 0;
    reg [260:0] temp50 = 0;
    reg [260:0] temp51 = 0;
    reg [260:0] temp52 = 0;
    reg [260:0] temp53 = 0;
    reg [260:0] temp54 = 0;
    reg [260:0] temp55 = 0;
    reg [260:0] temp56 = 0;
    reg [260:0] temp57 = 0;
    reg [260:0] temp58 = 0;
    reg [260:0] temp59 = 0;
    reg [260:0] temp60 = 0;
    reg [260:0] temp61 = 0;
    reg [260:0] temp62 = 0;
    reg [260:0] temp63 = 0;
    reg [260:0] temp64 = 0;
    reg [260:0] temp65 = 0;
    reg [260:0] temp66 = 0;
    reg [260:0] temp67 = 0;
    reg [260:0] temp68 = 0;
    reg [260:0] temp69 = 0;
    reg [260:0] temp70 = 0;
    reg [260:0] temp71 = 0;
    reg [260:0] temp72 = 0;
    reg [260:0] temp73 = 0;
    reg [260:0] temp74 = 0;


    
    reg [260:0] temp0_3 = 0;
    reg [260:0] temp4_7 = 0;
    reg [260:0] temp8_11 = 0;
    reg [260:0] temp12_15 = 0;
    reg [260:0] temp16_19 = 0;
    reg [260:0] temp20_23 = 0;
    reg [260:0] temp24_27 = 0;
    reg [260:0] temp28_31 = 0;
    reg [260:0] temp32_35 = 0;
    reg [260:0] temp36_39 = 0;
    reg [260:0] temp40_43 = 0;
    reg [260:0] temp44_47 = 0;
    reg [260:0] temp48_51 = 0;
    reg [260:0] temp52_55 = 0;
    reg [260:0] temp56_59 = 0;
    reg [260:0] temp60_63 = 0;
    reg [260:0] temp64_67 = 0;
    reg [260:0] temp68_71 = 0;
    reg [260:0] temp72_74 = 0;
    
    reg [260:0] temp0_15 = 0;
    reg [260:0] temp16_31 = 0;
    reg [260:0] temp32_47 = 0;
    reg [260:0] temp48_63 = 0;
    reg [260:0] temp64_74 = 0;
    reg [260:0] temp64_74_delay = 0;
    
    reg [260:0] temp0_63 = 0;
    
    reg [260:0] temp0_74 = 0;
    
    always@(posedge clk)
    begin
        if(reset == 1'b1)
        begin
            temp0 = 0;
            temp1 = 0;
            temp2 = 0;
            temp3 = 0;
            temp4 = 0;
            temp5 = 0;
            temp6 = 0;
            temp7 = 0;
            temp8 = 0;
            temp9 = 0;
            temp10 = 0;
            temp11 = 0;
            temp12 = 0;
            temp13 = 0;
            temp14 = 0;
            temp15 = 0;
            temp16 = 0;
            temp17 = 0;
            temp18 = 0;
            temp19 = 0;
            temp20 = 0;
            temp21 = 0;
            temp22 = 0;
            temp23 = 0;
            temp24 = 0;
            temp25 = 0;
            temp26 = 0;
            temp27 = 0;
            temp28 = 0;
            temp29 = 0;
            temp30 = 0;
            temp31 = 0;
            temp32 = 0;
            temp33 = 0;
            temp34 = 0;
            temp35 = 0;
            temp36 = 0;
            temp37 = 0;
            temp38 = 0;
            temp39 = 0;
            temp40 = 0;
            temp41 = 0;
            temp42 = 0;
            temp43 = 0;
            temp44 = 0;
            temp45 = 0;
            temp46 = 0;
            temp47 = 0;
            temp48 = 0;
            temp49 = 0;
            temp50 = 0;
            temp51 = 0;
            temp52 = 0;
            temp53 = 0;
            temp54 = 0;
            temp55 = 0;
            temp56 = 0;
            temp57 = 0;
            temp58 = 0;
            temp59 = 0;
            temp60 = 0;
            temp61 = 0;
            temp62 = 0;
            temp63 = 0;
            temp64 = 0;
            temp65 = 0;
            temp66 = 0;
            temp67 = 0;
            temp68 = 0;
            temp69 = 0;
            temp70 = 0;
            temp71 = 0;
            temp72 = 0;
            temp73 = 0;
            temp74 = 0;
            temp0_3 = 0;
            temp4_7 = 0;
            temp8_11 = 0;
            temp12_15 = 0;
            temp16_19 = 0;
            temp20_23 = 0;
            temp24_27 = 0;
            temp28_31 = 0;
            temp32_35 = 0;
            temp36_39 = 0;
            temp40_43 = 0;
            temp44_47 = 0;
            temp48_51 = 0;
            temp52_55 = 0;
            temp56_59 = 0;
            temp60_63 = 0;
            temp64_67 = 0;
            temp68_71 = 0;
            temp72_74 = 0;
            temp0_15 = 0;
            temp16_31 = 0;
            temp32_47 = 0;
            temp48_63 = 0;
            temp64_74 = 0;
            temp0_63 = 0;
            temp0_74 = 0;
            temp64_74_delay = 0;
        end
        
        else   
        begin
            temp0 <= ((x[0])?x0:0)+ ((x[1])?x1:0)+ ((x[2])?x2:0)+ ((x[3])?x3:0); 
            temp1 <= ((x[4])?x4:0)+ ((x[5])?x5:0)+ ((x[6])?x6:0)+ ((x[7])?x7:0); 
            temp2 <= ((x[8])?x8:0)+ ((x[9])?x9:0)+ ((x[10])?x10:0)+ ((x[11])?x11:0); 
            temp3 <= ((x[12])?x12:0)+ ((x[13])?x13:0)+ ((x[14])?x14:0)+ ((x[15])?x15:0); 
            temp4 <= ((x[16])?x16:0)+ ((x[17])?x17:0)+ ((x[18])?x18:0)+ ((x[19])?x19:0); 
            temp5 <= ((x[20])?x20:0)+ ((x[21])?x21:0)+ ((x[22])?x22:0)+ ((x[23])?x23:0); 
            temp6 <= ((x[24])?x24:0)+ ((x[25])?x25:0)+ ((x[26])?x26:0)+ ((x[27])?x27:0); 
            temp7 <= ((x[28])?x28:0)+ ((x[29])?x29:0)+ ((x[30])?x30:0)+ ((x[31])?x31:0); 
            temp8 <= ((x[32])?x32:0)+ ((x[33])?x33:0)+ ((x[34])?x34:0)+ ((x[35])?x35:0); 
            temp9 <= ((x[36])?x36:0)+ ((x[37])?x37:0)+ ((x[38])?x38:0)+ ((x[39])?x39:0); 
            temp10 <= ((x[40])?x40:0)+ ((x[41])?x41:0)+ ((x[42])?x42:0)+ ((x[43])?x43:0); 
            temp11 <= ((x[44])?x44:0)+ ((x[45])?x45:0)+ ((x[46])?x46:0)+ ((x[47])?x47:0); 
            temp12 <= ((x[48])?x48:0)+ ((x[49])?x49:0)+ ((x[50])?x50:0)+ ((x[51])?x51:0); 
            temp13 <= ((x[52])?x52:0)+ ((x[53])?x53:0)+ ((x[54])?x54:0)+ ((x[55])?x55:0); 
            temp14 <= ((x[56])?x56:0)+ ((x[57])?x57:0)+ ((x[58])?x58:0)+ ((x[59])?x59:0); 
            temp15 <= ((x[60])?x60:0)+ ((x[61])?x61:0)+ ((x[62])?x62:0)+ ((x[63])?x63:0); 
            temp16 <= ((x[64])?x64:0)+ ((x[65])?x65:0)+ ((x[66])?x66:0)+ ((x[67])?x67:0); 
            temp17 <= ((x[68])?x68:0)+ ((x[69])?x69:0)+ ((x[70])?x70:0)+ ((x[71])?x71:0); 
            temp18 <= ((x[72])?x72:0)+ ((x[73])?x73:0)+ ((x[74])?x74:0)+ ((x[75])?x75:0); 
            temp19 <= ((x[76])?x76:0)+ ((x[77])?x77:0)+ ((x[78])?x78:0)+ ((x[79])?x79:0); 
            temp20 <= ((x[80])?x80:0)+ ((x[81])?x81:0)+ ((x[82])?x82:0)+ ((x[83])?x83:0); 
            temp21 <= ((x[84])?x84:0)+ ((x[85])?x85:0)+ ((x[86])?x86:0)+ ((x[87])?x87:0); 
            temp22 <= ((x[88])?x88:0)+ ((x[89])?x89:0)+ ((x[90])?x90:0)+ ((x[91])?x91:0); 
            temp23 <= ((x[92])?x92:0)+ ((x[93])?x93:0)+ ((x[94])?x94:0)+ ((x[95])?x95:0); 
            temp24 <= ((x[96])?x96:0)+ ((x[97])?x97:0)+ ((x[98])?x98:0)+ ((x[99])?x99:0); 
            temp25 <= ((x[100])?x100:0)+ ((x[101])?x101:0)+ ((x[102])?x102:0)+ ((x[103])?x103:0); 
            temp26 <= ((x[104])?x104:0)+ ((x[105])?x105:0)+ ((x[106])?x106:0)+ ((x[107])?x107:0); 
            temp27 <= ((x[108])?x108:0)+ ((x[109])?x109:0)+ ((x[110])?x110:0)+ ((x[111])?x111:0); 
            temp28 <= ((x[112])?x112:0)+ ((x[113])?x113:0)+ ((x[114])?x114:0)+ ((x[115])?x115:0); 
            temp29 <= ((x[116])?x116:0)+ ((x[117])?x117:0)+ ((x[118])?x118:0)+ ((x[119])?x119:0); 
            temp30 <= ((x[120])?x120:0)+ ((x[121])?x121:0)+ ((x[122])?x122:0)+ ((x[123])?x123:0); 
            temp31 <= ((x[124])?x124:0)+ ((x[125])?x125:0)+ ((x[126])?x126:0)+ ((x[127])?x127:0); 
            temp32 <= ((x[128])?x128:0)+ ((x[129])?x129:0)+ ((x[130])?x130:0)+ ((x[131])?x131:0); 
            temp33 <= ((x[132])?x132:0)+ ((x[133])?x133:0)+ ((x[134])?x134:0)+ ((x[135])?x135:0); 
            temp34 <= ((x[136])?x136:0)+ ((x[137])?x137:0)+ ((x[138])?x138:0)+ ((x[139])?x139:0); 
            temp35 <= ((x[140])?x140:0)+ ((x[141])?x141:0)+ ((x[142])?x142:0)+ ((x[143])?x143:0); 
            temp36 <= ((x[144])?x144:0)+ ((x[145])?x145:0)+ ((x[146])?x146:0)+ ((x[147])?x147:0); 
            temp37 <= ((x[148])?x148:0)+ ((x[149])?x149:0)+ ((x[150])?x150:0)+ ((x[151])?x151:0); 
            temp38 <= ((x[152])?x152:0)+ ((x[153])?x153:0)+ ((x[154])?x154:0)+ ((x[155])?x155:0); 
            temp39 <= ((x[156])?x156:0)+ ((x[157])?x157:0)+ ((x[158])?x158:0)+ ((x[159])?x159:0); 
            temp40 <= ((x[160])?x160:0)+ ((x[161])?x161:0)+ ((x[162])?x162:0)+ ((x[163])?x163:0); 
            temp41 <= ((x[164])?x164:0)+ ((x[165])?x165:0)+ ((x[166])?x166:0)+ ((x[167])?x167:0); 
            temp42 <= ((x[168])?x168:0)+ ((x[169])?x169:0)+ ((x[170])?x170:0)+ ((x[171])?x171:0); 
            temp43 <= ((x[172])?x172:0)+ ((x[173])?x173:0)+ ((x[174])?x174:0)+ ((x[175])?x175:0); 
            temp44 <= ((x[176])?x176:0)+ ((x[177])?x177:0)+ ((x[178])?x178:0)+ ((x[179])?x179:0); 
            temp45 <= ((x[180])?x180:0)+ ((x[181])?x181:0)+ ((x[182])?x182:0)+ ((x[183])?x183:0); 
            temp46 <= ((x[184])?x184:0)+ ((x[185])?x185:0)+ ((x[186])?x186:0)+ ((x[187])?x187:0); 
            temp47 <= ((x[188])?x188:0)+ ((x[189])?x189:0)+ ((x[190])?x190:0)+ ((x[191])?x191:0); 
            temp48 <= ((x[192])?x192:0)+ ((x[193])?x193:0)+ ((x[194])?x194:0)+ ((x[195])?x195:0); 
            temp49 <= ((x[196])?x196:0)+ ((x[197])?x197:0)+ ((x[198])?x198:0)+ ((x[199])?x199:0); 
            temp50 <= ((x[200])?x200:0)+ ((x[201])?x201:0)+ ((x[202])?x202:0)+ ((x[203])?x203:0); 
            temp51 <= ((x[204])?x204:0)+ ((x[205])?x205:0)+ ((x[206])?x206:0)+ ((x[207])?x207:0); 
            temp52 <= ((x[208])?x208:0)+ ((x[209])?x209:0)+ ((x[210])?x210:0)+ ((x[211])?x211:0); 
            temp53 <= ((x[212])?x212:0)+ ((x[213])?x213:0)+ ((x[214])?x214:0)+ ((x[215])?x215:0); 
            temp54 <= ((x[216])?x216:0)+ ((x[217])?x217:0)+ ((x[218])?x218:0)+ ((x[219])?x219:0); 
            temp55 <= ((x[220])?x220:0)+ ((x[221])?x221:0)+ ((x[222])?x222:0)+ ((x[223])?x223:0); 
            temp56 <= ((x[224])?x224:0)+ ((x[225])?x225:0)+ ((x[226])?x226:0)+ ((x[227])?x227:0); 
            temp57 <= ((x[228])?x228:0)+ ((x[229])?x229:0)+ ((x[230])?x230:0)+ ((x[231])?x231:0); 
            temp58 <= ((x[232])?x232:0)+ ((x[233])?x233:0)+ ((x[234])?x234:0)+ ((x[235])?x235:0); 
            temp59 <= ((x[236])?x236:0)+ ((x[237])?x237:0)+ ((x[238])?x238:0)+ ((x[239])?x239:0); 
            temp60 <= ((x[240])?x240:0)+ ((x[241])?x241:0)+ ((x[242])?x242:0)+ ((x[243])?x243:0); 
            temp61 <= ((x[244])?x244:0)+ ((x[245])?x245:0)+ ((x[246])?x246:0)+ ((x[247])?x247:0); 
            temp62 <= ((x[248])?x248:0)+ ((x[249])?x249:0)+ ((x[250])?x250:0)+ ((x[251])?x251:0); 
            temp63 <= ((x[252])?x252:0)+ ((x[253])?x253:0)+ ((x[254])?x254:0)+ ((x[255])?x255:0); 
            temp64 <= ((x[256])?x256:0)+ ((x[257])?x257:0)+ ((x[258])?x258:0)+ ((x[259])?x259:0); 
            temp65 <= ((x[260])?x260:0)+ ((x[261])?x261:0)+ ((x[262])?x262:0)+ ((x[263])?x263:0); 
            temp66 <= ((x[264])?x264:0)+ ((x[265])?x265:0)+ ((x[266])?x266:0)+ ((x[267])?x267:0); 
            temp67 <= ((x[268])?x268:0)+ ((x[269])?x269:0)+ ((x[270])?x270:0)+ ((x[271])?x271:0); 
            temp68 <= ((x[272])?x272:0)+ ((x[273])?x273:0)+ ((x[274])?x274:0)+ ((x[275])?x275:0); 
            temp69 <= ((x[276])?x276:0)+ ((x[277])?x277:0)+ ((x[278])?x278:0)+ ((x[279])?x279:0); 
            temp70 <= ((x[280])?x280:0)+ ((x[281])?x281:0)+ ((x[282])?x282:0)+ ((x[283])?x283:0); 
            temp71 <= ((x[284])?x284:0)+ ((x[285])?x285:0)+ ((x[286])?x286:0)+ ((x[287])?x287:0); 
            temp72 <= ((x[288])?x288:0)+ ((x[289])?x289:0)+ ((x[290])?x290:0)+ ((x[291])?x291:0); 
            temp73 <= ((x[292])?x292:0)+ ((x[293])?x293:0)+ ((x[294])?x294:0)+ ((x[295])?x295:0); 
            temp74 <= ((x[296])?x296:0)+ ((x[297])?x297:0)+ ((x[298])?x298:0)+ ((x[299])?x299:0);  
                   
            temp0_3 <= temp0 + temp1 + temp2 + temp3;
            temp4_7 <= temp4 + temp5 + temp6 + temp7;
            temp8_11 <= temp8 + temp9 + temp10 + temp11;
            temp12_15 <= temp12 + temp13 + temp14 + temp15;
            temp16_19 <= temp16 + temp17 + temp18 + temp19;
            temp20_23 <= temp20 + temp21 + temp22 + temp23;
            temp24_27 <= temp24 + temp25 + temp26 + temp27;
            temp28_31 <= temp28 + temp29 + temp30 + temp31;
            temp32_35 <= temp32 + temp33 + temp34 + temp35;
            temp36_39 <= temp36 + temp37 + temp38 + temp39;
            temp40_43 <= temp40 + temp41 + temp42 + temp43;
            temp44_47 <= temp44 + temp45 + temp46 + temp47;
            temp48_51 <= temp48 + temp49 + temp50 + temp51;
            temp52_55 <= temp52 + temp53 + temp54 + temp55;
            temp56_59 <= temp56 + temp57 + temp58 + temp59;
            temp60_63 <= temp60 + temp61 + temp62 + temp63;
            temp64_67 <= temp64 + temp65 + temp66 + temp67;
            temp68_71 <= temp68 + temp69 + temp70 + temp71;
            temp72_74 <= temp72 + temp73 + temp74;
            
            temp0_15 <= temp0_3 + temp4_7 + temp8_11 + temp12_15;
            temp16_31 <= temp16_19 + temp20_23 + temp24_27 + temp28_31;
            temp32_47 <= temp32_35 + temp36_39 + temp40_43 + temp44_47;
            temp48_63 <= temp48_51 + temp52_55 + temp56_59 + temp60_63;
            temp64_74 <= temp64_67 + temp68_71 + temp72_74;
            temp64_74_delay <= temp64_74;
            //Delay by 1 CLK cycle, since we need to synchronise the temp0_63 and temp64_74
    
            temp0_63 <= temp0_15 + temp16_31 + temp32_47 + temp48_63;
            temp0_74 <= temp0_63 + temp64_74_delay;
       end 
    end
    
    assign o = temp0_74;
endmodule
